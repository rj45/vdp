// from: https://github.com/lawrie/ulx3s_zx_spectrum/
// Original origin / license unknown

`default_nettype none
`timescale 1ns / 1ps

// module port
//
module hdmi(
  input  logic clk_pix,
  input  logic clk_pix5x,
  input  logic rst_pix,
  input  logic rst_pix5x,
  input  logic [7:0] r, g, b,
  input  logic de, hsync, vsync,
  output logic [3:0] gpdi_dp, gpdi_dn
);

    logic [7:0] r_r;
    logic [7:0] g_r;
    logic [7:0] b_r;
    logic       de_r;
    logic       hsync_r;
    logic       vsync_r;

    // register inputs to improve performance
    always_ff @(posedge clk_pix) begin
        r_r     <= r;
        g_r     <= g;
        b_r     <= b;
        de_r    <= de;
        hsync_r <= hsync;
        vsync_r <= vsync;
    end

    // 10b8b TMDS encoding of RGB and Sync
    //
    wire [9:0] TMDS_red, TMDS_green, TMDS_blue;
    tmds_encoder encode_R(.clk(clk_pix), .i_reset(rst_pix), .VD(r_r), .CD(2'b00)            , .VDE(de_r), .TMDS(TMDS_red));
    tmds_encoder encode_G(.clk(clk_pix), .i_reset(rst_pix), .VD(g_r), .CD(2'b00)            , .VDE(de_r), .TMDS(TMDS_green));
    tmds_encoder encode_B(.clk(clk_pix), .i_reset(rst_pix), .VD(b_r), .CD({vsync_r,hsync_r}), .VDE(de_r), .TMDS(TMDS_blue));

    smoldvi_clock_driver ser_ck (
    	.clk_x5    (clk_pix5x),
    	.rst_n_x5  (~rst_pix5x),

    	.qp        (gpdi_dp[3]),
    	.qn        (gpdi_dn[3])
    );

    smoldvi_serialiser ser_red (
    	.clk_pix   (clk_pix),
    	.rst_n_pix (~rst_pix),
    	.clk_x5    (clk_pix5x),
    	.rst_n_x5  (~rst_pix5x),

    	.d         (TMDS_red),
    	.qp        (gpdi_dp[2]),
    	.qn        (gpdi_dn[2])
    );

    smoldvi_serialiser ser_green (
    	.clk_pix   (clk_pix),
    	.rst_n_pix (~rst_pix),
    	.clk_x5    (clk_pix5x),
    	.rst_n_x5  (~rst_pix5x),

    	.d         (TMDS_green),
    	.qp        (gpdi_dp[1]),
    	.qn        (gpdi_dn[1])
    );

    smoldvi_serialiser ser_blue (
    	.clk_pix   (clk_pix),
    	.rst_n_pix (~rst_pix),
    	.clk_x5    (clk_pix5x),
    	.rst_n_x5  (~rst_pix5x),

    	.d         (TMDS_blue),
    	.qp        (gpdi_dp[0]),
    	.qn        (gpdi_dn[0])
    );

endmodule

// tmds_encoder performs Transition-minimized differential signaling (TMDS) encoding of
// 8-bits of pixel data and 2-bits of control data to a 10-bit TMDS encoded format.
// Requires synthesizing with System Verilog 2017.
// (this module is unit tested with cocotb framework)
//
// Borrowed from: https://github.com/juj/gowin_flipflop_drainer/blob/main/src/hdmi.v#L1-L221
// License:
//   All code in this repository is released to public domain. Do with it whatever you wish. No attributions.
module tmds_encoder(
  input clk,         // HDMI pixel clock
  input i_reset,            // reset (active high)
  input [7:0] VD,       // Input 8-bit color
  input [1:0] CD,       // control data (vsync and hsync)
  input VDE,   // high=pixel data active. low=display is in blanking area
  output reg [9:0] TMDS   // encoded 10-bit TMDS data
);
  // Intermediate pipelined variables: the number after each reg specifies the clock cycle of the pipeline the values are accessed at.

  // Reset
  reg rst0;
  // Unencoded input data
  reg [7:0] dat0, dat1, dat2, dat3, dat4, dat5, dat6, dat7 ;
  // Control signal (hsync and vsync)
  reg [1:0] ctl0, ctl1, ctl2, ctl3, ctl4, ctl5, ctl6, ctl7, ctl8, ctl9, ctl10, ctl11, ctl12, ctl13, ctl14, ctl15, ctl16, ctl17, ctl18;
  // Display enable signal
  reg den0, den1, den2, den3, den4, den5, den6, den7, den8, den9, den10, den11, den12, den13, den14, den15, den16, den17, not_den18;
  // Parity count of input data
  reg [4:0] par1, par2, par3, par4, par5, par6, par7, par8;
  // Parity bit of input data (if set, input had >= 4 bits set).
  reg par9, par10, par11, par12, par13, par14, par15, par16, par17, par18;
  // Intermediate encoded stage of the input vector.
  reg [7:0] enc3, enc4, enc5, enc6, enc7, enc8, enc9, enc10, enc11, enc12, enc13, enc14, enc15, enc16, enc17, enc18;
  // Count the number of ones in the intermediate encoded data
  reg signed [3:0] eon10, eon11, eon13, eon14, eon15, eon16, eon17, eon18;
  // Is Encoded ONes even?
  reg eve18;
  // Temp values for accumulating the count of ones in the encoded vector.
  reg [3:0] tpa10, tpa11, tpb11;
  reg [2:0] tpa12, tpb12;
  // Pipelined values for updating the bias count.
  reg signed [3:0] inv18, shr18, shl18;
  // Pipelined values for the output TMDS data.
  reg [9:0] tmds_blank18, tmds_even18, tmds_pos18, tmds_neg18;
  // 'bias' stores the running TMDS ones vs zeros balance count. If > 0, we've sent more ones to the bus,
  // if < 0, we've sent more zeroes than ones, if == 0, we are at equal balance.
  reg signed [3:0] bias;

  always_ff @(posedge clk) begin
    // Clock 0: register inputs
    rst0 <= i_reset;
    dat0 <= VD;
    ctl0 <= CD;
    den0 <= VDE;

    // Clock 1: handle reset early by folding it into the other fields
    dat1 <= dat0;
    ctl1 <= rst0 ? 2'b0 : ctl0;
    den1 <= rst0 ? 1'b0 : den0;

    // Clock 2: sanitize image data to zero if inside display blank (or reset)
    dat2 <= den1 ? dat1 : 8'b0;
    ctl2 <= ctl1;
    den2 <= den1;

    // Clocks 3-7: Pipeline 'dat' for the duration of the parity encoding below.
    dat3 <= dat2;
    dat4 <= dat3;
    dat5 <= dat4;
    dat6 <= dat5;
    dat7 <= dat6;

    // Clocks 1-8: Calculate parity, i.e. whether the input vector 'dat' has more
    //             ones in it than zeros. If it has 4 zeros and 4 ones, use ~dat[0]
    //             as a tie. To do that, start with constant vector 00001, and for
    //             each bit set in input 'dat', shift 'par' left by one place, filling
    //             in ones. At the end par[4] will specifies whether there were more
    //             ones than zeroes.
    par1 <= 5'b00001;
    par2 <= dat1[1] ? {par1[3:0], 1'b1} : par1; // = 000ab (a,b=unknown, 000=zeroes)
    par3 <= dat2[2] ? {par2[3:0], 1'b1} : par2; // = 00abc
    par4 <= dat3[3] ? {par3[3:0], 1'b1} : par3; // = 0abcd
    par5 <= dat4[4] ? {par4[3:0], 1'b1} : par4; // = abcdx (x=don't care, rely on optimizer to clear these away)
    par6 <= dat5[5] ? {par5[3:0], 1'b1} : par5; // = bcdxx
    par7 <= dat6[6] ? {par6[3:0], 1'b1} : par6; // = cdxxx
    par8 <= dat7[7] ? {par7[3:0], 1'b1} : par7; // = dxxxx

    // Clocks 9-18: No further calculation needed for parity. Keep pipelining it forward
    //              in a single bit vector.
    par9 <= par8[4]; // At the end of computation par[4] records the parity.
    par10 <= par9;
    par11 <= par10;
    par12 <= par11;
    par13 <= par12;
    par14 <= par13;
    par15 <= par14;
    par16 <= par15;
    par17 <= par16;
    par18 <= par17;

    // Clocks 3-18: No more changes needed to the Display Enable signal, flow it through the pipeline
    den3 <= den2;
    den4 <= den3;
    den5 <= den4;
    den6 <= den5;
    den7 <= den6;
    den8 <= den7;
    den9 <= den8;
    den10 <= den9;
    den11 <= den10;
    den12 <= den11;
    den13 <= den12;
    den14 <= den13;
    den15 <= den14;
    den16 <= den15;
    den17 <= den16;
    not_den18 <= ~den17;

    // Clocks 3-18: Pipeline ctrl data (hsync & vsync), no changes needed.
    ctl3 <= ctl2;
    ctl4 <= ctl3;
    ctl5 <= ctl4;
    ctl6 <= ctl5;
    ctl7 <= ctl6;
    ctl8 <= ctl7;
    ctl9 <= ctl8;
    ctl10 <= ctl9;
    ctl11 <= ctl10;
    ctl12 <= ctl11;
    ctl13 <= ctl12;
    ctl14 <= ctl13;
    ctl15 <= ctl14;
    ctl16 <= ctl15;
    ctl17 <= ctl16;
    ctl18 <= ctl17;

    // Clocks 3-9: perform intermediate encoded vector 'enc' of the input 'data' field. At the
    //             end of the encoding, the DVI spec says the encoded vector should look like
    //             follows:
    // enc <= { parity ^ data[0] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[7],
    //                   data[0] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[6],
    //          parity ^ data[0] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[5],
    //                   data[0] ^ data[1] ^ data[2] ^ data[3] ^ data[4],
    //          parity ^ data[0] ^ data[1] ^ data[2] ^ data[3],
    //                   data[0] ^ data[1] ^ data[2],
    //          parity ^ data[0] ^ data[1],
    //                   data[0] };
    //
    // Calculate it across a few clock cycles to avoid high complexity per clock. (ignore parity first)
    // Bit lanes after each clock cycle:
    //                [7]     [6]    [5]   [4]  [3] [2] [1] [0]
    // Clock 2:        7       6      5     4    3   2   1   0
    // Clock 3:       76      65     54    43   32  21  10   0
    // Clock 4:     7654    6543   5432  4321 3210 210  10   0
    // Clock 5: 76543210 6543210 543210 43210 3210 210  10   0

    enc3 <= {dat2[7:1]^dat2[6:0], dat2[  0]};
    enc4 <= {enc3[7:2]^enc3[5:0], enc3[1:0]};
    enc5 <= {enc4[7:4]^enc4[3:0], enc4[3:0]};
    enc6 <= enc5;
    enc7 <= enc6;
    enc8 <= enc7;

    // Clock 9: Meanwhile, parity computation has completed, so apply the final parity XOR to the
    //          intermediate encoded vector.
    enc9 <= enc8 ^ {4{par8[4], 1'b0}};
    enc10 <= enc9;
    enc11 <= enc10;
    enc12 <= enc11;
    enc13 <= enc12;
    enc14 <= enc13;
    enc15 <= enc14;
    enc16 <= enc15;
    enc17 <= enc16;
    enc18 <= enc17;

    // Clocks 10-17: calculate 'eon' (Encoded ONes vs zeros): a signed count that specifies whether
    //               vector 'enc' has more ones or zeroes in it.
    tpa10 <= enc9[3:0] ^ enc9[7:4]; // Fold the 8 bit enc vector into two 4-bit halves, and half-
    tpa11 <= tpa10;     // Then calculate the number of ones in them in parallel
    tpb11 <= enc10[3:0] & enc10[7:4];//tpb10;
    tpa12 <= $countones(tpa11);     // Then calculate the number of ones in them in parallel
    tpb12 <= $countones(tpb11);
    eon13 <= tpa12 + {tpb12, 1'b0}; // Then use a 3-bit + 4-bit addition to bring the full count.
    eon14 <= eon13 - 3'd4;          // And make the result signed.
    eon15 <= eon14;
    eon16 <= eon15;
    eon17 <= eon16;
    eon18 <= eon17;

    // 'eon17' is a count of balance of ones vs zeros in input encoded vector 'enc':
    //        #ones: 8 7 6 5 4  3  2  1  0
    // #ones-#zeros: 8 6 4 2 0 -2 -4 -6 -8
    // value of eon: 4 3 2 1 0 -1 -2 -3 -4

    // Pipeline a few finishing touches:
    eve18 <= eon17 == 0;                      // is the balance equal (zero)?
    inv18 <= par17 ? -eon17     : eon17;      // invert balance count based on parity.
    shr18 <= par17 ? eon17      : eon17-1'b1; // right shift balance count based on parity.
    shl18 <= par17 ? eon17-1'b1 : eon17;      // left shift balance count based on parity.
    tmds_blank18 <= {~ctl17[1], 9'b101010100} ^ {10{ctl17[0]}};
    tmds_even18 <= {par17, ~par17, {8{par17}} ^ enc17};
    tmds_pos18 <= {1'b1, ~par17, 8'hff ^ enc17};
    tmds_neg18 <= {1'b0, ~par17,         enc17};

    // Clocks 14-17 above:
    // These are "empty" filler clock stages that contain no computations on any of the variables,
    // but they only perform direct passthrough of the values that have been computed so far.
    // Gowin IDE Analyzer reports that this improves max. timing performance.

    // Clock 18: finally output the TMDS encoded value, and update bias value
    if (not_den18) begin // In display blank?
      TMDS <= tmds_blank18;              // Output control words for hsync and vsync
      bias <= 0;                           // Bias resets to zero in blank
    end else if (eve18 || bias == 0) begin // If current bias is even, or encoded balance is even..
      TMDS <= tmds_even18;               // .. use a specific 'even' state TMDS formula.
      bias <= bias + inv18;                // This does not seem to be strictly necessary, you can try removing this else block for tiny bit more performance.
    end else if (bias[3] == eon18[3]) begin // Otherwise, noneven bias and balance, so use the main TMDS encoding formula
      TMDS <= tmds_pos18;
      bias <= bias - shr18; // and update running bias of ones vs zeros sent.
    end else begin
      TMDS <= tmds_neg18;
      bias <= bias + shl18;
    end
  end
endmodule



//--------------------------------------------------------------------------------
// Engineer: Mike Field <hamster@snap.net.nz>
//
// Description: TMDS Encoder
//     8 bits colour, 2 control bits and one blanking bits in
//       10 bits of TMDS encoded data out
//     Clocked at the pixel clock
//
//--------------------------------------------------------------------------------
// See: http://hamsterworks.co.nz/mediawiki/index.php/Dvid_test
//      http://hamsterworks.co.nz/mediawiki/index.php/FPGA_Projects
//
// Copyright (c) 2012 Mike Field <hamster@snap.net.nz>
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.

// module tmds_encoder(
//     input  logic clk,
//     input  logic i_reset,
//     input  logic [7:0] VD,
//     input  logic [1:0] CD,
//     input  logic VDE,
//     output logic [9:0] TMDS
// );
//     logic [8:0] xored;
//     logic [8:0] xnored;
//     logic [3:0] ones;
//     logic [8:0] data_word;
//     logic [8:0] data_word_inv;
//     logic [3:0] data_word_disparity;
//     logic [3:0] dc_bias = 1'b0;

//     // Work out the two different encodings for the byte
//     assign xored[0] = VD[0];
//     assign xored[1] = VD[1] ^ xored[0];
//     assign xored[2] = VD[2] ^ xored[1];
//     assign xored[3] = VD[3] ^ xored[2];
//     assign xored[4] = VD[4] ^ xored[3];
//     assign xored[5] = VD[5] ^ xored[4];
//     assign xored[6] = VD[6] ^ xored[5];
//     assign xored[7] = VD[7] ^ xored[6];
//     assign xored[8] = 1'b1;
//     assign xnored[0] = VD[0];
//     assign xnored[1] = ~(VD[1] ^ xnored[0]);
//     assign xnored[2] = ~(VD[2] ^ xnored[1]);
//     assign xnored[3] = ~(VD[3] ^ xnored[2]);
//     assign xnored[4] = ~(VD[4] ^ xnored[3]);
//     assign xnored[5] = ~(VD[5] ^ xnored[4]);
//     assign xnored[6] = ~(VD[6] ^ xnored[5]);
//     assign xnored[7] = ~(VD[7] ^ xnored[6]);
//     assign xnored[8] = 1'b0;
//     // Count how many ones are set in data
//     assign ones = 4'b0000 +
//         VD[0] + VD[1] + VD[2] + VD[3] +
//         VD[4] + VD[5] + VD[6] + VD[7];
//     // Decide which encoding to use
//     always @(ones, VD[0], xnored, xored) begin
//     if (ones > 4 || (ones == 4 && VD[0] == 1'b0)) begin
//         data_word <= xnored;
//         data_word_inv <=  ~(xnored);
//     end
//     else begin
//         data_word <= xored;
//         data_word_inv <=  ~(xored);
//     end
//     end

//     // Work out the DC bias of the dataword;
//     assign data_word_disparity = 4'b1100 +
//         data_word[0] + data_word[1] + data_word[2] + data_word[3] +
//         data_word[4] + data_word[5] + data_word[6] + data_word[7];
//     // Now work out what the output should be
//     always @(posedge clk) begin
//         if (VDE == 1'b0) begin
//             // In the control periods, all values have and have balanced bit count
//             case(CD)
//                 2'b00 : begin
//                     TMDS <= 10'b1101010100;
//                 end
//                 2'b01 : begin
//                     TMDS <= 10'b0010101011;
//                 end
//                 2'b10 : begin
//                     TMDS <= 10'b0101010100;
//                 end
//                 default : begin
//                     TMDS <= 10'b1010101011;
//                 end
//             endcase
//             dc_bias <= {4{1'b0}};
//         end else begin
//             if (dc_bias == 5'b00000 || data_word_disparity == 0) begin
//                 // dataword has no disparity
//                 if (data_word[8] == 1'b1) begin
//                     TMDS <= {2'b01,data_word[7:0]};
//                     dc_bias <= dc_bias + data_word_disparity;
//                 end else begin
//                     TMDS <= {2'b10,data_word_inv[7:0]};
//                     dc_bias <= dc_bias - data_word_disparity;
//                 end
//             end else if (
//                 (dc_bias[3] == 1'b0 && data_word_disparity[3] == 1'b0) ||
//                 (dc_bias[3] == 1'b1 && data_word_disparity[3] == 1'b1)
//             ) begin
//                 TMDS <= {1'b1,data_word[8],data_word_inv[7:0]};
//                 dc_bias <= dc_bias + data_word[8] - data_word_disparity;
//             end else begin
//                 TMDS <= {1'b0,data_word};
//                 dc_bias <= dc_bias - data_word_inv[8] + data_word_disparity;
//             end
//         end
//     end
// endmodule
